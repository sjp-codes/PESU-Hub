module gate(y,a,b);
input a,b;
output y;
assign y = -------;
endmodule